module HitDetection_updated (
    input clk,

    input [9:0] x1, // of top left corner 
    input [9:0] x2,

	
    input p1_attack_flag,
    input p2_attack_flag,
		 
    input p1_dir_attack,
    input p2_dir_attack,
	 
	 // must input state to check if player is blocking or under recovery
	 // if its easier to get the respective flags corresponding to these states then lemme know or you can
	 // change the code appropriately I made it so it can be easily changed. Its very dynamically written so its super cool
	 
	 //combined input:
	 input [3:0] state1,
	 input [3:0] state2,

    output reg [1:0] p1_stunmode,
    output reg [1:0] p2_stunmode

);

    localparam 
		SCREEN_WIDTH 			= 10'd640,
		SCREEN_HEIGHT        = 10'd480,

		neutral_HITBOX_WIDTH = 10'd30,
    	dir_HITBOX_WIDTH     = 10'd48,
    	HITBOX_HEIGHT        = 10'd80,

    	BASE_WIDTH           = 10'd64, 
    	PLAYER_HEIGHT        = 10'd240,

		S_BACKWARD           = 4'd2,
		S_Attack_recovery    = 4'd5;


	// stunmode: 00 = neutral, 01 = hitstun, 10 = blockstun, 11 = whiff
	// if player is in whiff mode their hurtbox becomes the combined neutral hurt box and the attack_hitbox
	// i dont really need to indicate whiff mode but its there just in case we need it

	wire p1_blocking, p2_blocking;
	wire [1:0] attack_case;
	wire [9:0] attack_width, p1Hrtbox, p2Hrtbox;
	
	assign attack_case = {(p2_dir_attack | p2_attack_flag), (p1_dir_attack | p1_attack_flag)};
	assign attack_width = (p2_dir_attack | p1_dir_attack) ? dir_HITBOX_WIDTH : neutral_HITBOX_WIDTH;
	assign p1_blocking = state1 == S_BACKWARD;
	assign p2_blocking = state2 == S_BACKWARD;
//	assign p1_recov = state1 == S_Attack_recovery;
//	assign p2_recov = state2 == S_Attack_recovery;
	
	assign p1Hrtbox = (state1 == S_Attack_recovery) ? x1 + BASE_WIDTH + attack_width : x1 + BASE_WIDTH;
	assign p2Hrtbox = (state2 == S_Attack_recovery) ? x2 - attack_width : x2;


	initial begin
		p1_stunmode          = 2'b00;
		p2_stunmode          = 2'b00;
	end

	
	always @(posedge clk) begin	
		
		case(attack_case)
			
			2'b01: begin // p1 attack
				// check if p2 is within p1's attack hitbox
				if (x1 + BASE_WIDTH + attack_width > p2Hrtbox) begin
					if (~p2_blocking) begin 
						p1_stunmode = 2'b00; // p1's attack connnected
						p2_stunmode = 2'b01; // p2 in hitstun
						
					end else begin
						p1_stunmode = 2'b00; // p1's attack connnected
						p2_stunmode = 2'b10; // p2 in blockstun
					end
				end
			end
			
			2'b10: begin //p2 attack
				if (x2 - attack_width < p1Hrtbox) begin // attack connected
						if (~p1_blocking) begin 
							p2_stunmode = 2'b11; // atk connected
							p1_stunmode = 2'b01; // p1 in hitsun
						end else begin
							p2_stunmode = 2'b11; // p2's atk connnected
							p1_stunmode = 2'b10; // p2 in blockstun
						end
					end
			end
			
			2'b11: begin // both attacking simultaneously
				if (x1 + BASE_WIDTH + attack_width > x2 - attack_width) begin 
					// in this case both attacks connect and both players get damage
					p1_stunmode = 2'b01;
					p2_stunmode = 2'b01;
				end
			end	
			default: begin 
				p1_stunmode = 2'b00;
				p2_stunmode = 2'b00;
			end
		endcase
	end
		
endmodule
